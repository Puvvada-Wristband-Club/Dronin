/*
This is the NODE module for our network that handles the computations for each 
node. The PE(s) and IF module(s) are located here.
*/
`include "connect_parameters.v"


module node_module(N_clk, N_rst, if_i_flit, 
					if_i_credit, if_o_credit_valid,
					if_o_credit, if_o_data, if_o_data_valid, Node_id,
					a_in, a_out, dummy);
	
	localparam vc_bits = (`NUM_VCS > 1) ? $clog2(`NUM_VCS) : 1;
	  reg [vc_bits-1:0]   vc;


	input wire N_clk, N_rst;
	input wire [72:0] if_i_flit;
	input wire [7:0] Node_id;
	input wire [63:0] a_in;

	output wire [2:0] if_i_credit;
	output wire if_o_credit_valid;
	output wire [2:0] if_o_credit;
	output wire [72:0] if_o_data;
	output wire if_o_data_valid;
	output [63:0] a_out;
	output reg [63:0] dummy;
	
	reg [31:0] test_value_A = 32'b01000000001000000000000000000000; 
	reg [31:0] test_value_B = 32'b01000000100000000000000000000000;
	reg [31:0] test_value_C = 32'b00111111100100000000000000000000;
	
	// Local values for computation
	reg [63:0] a;
	assign a_out = a;

	wire req_ack;
	wire [31:0] PE_mult_result, PE_add_result;
	reg [31:0] send_data;
	reg [3:0] flit_count;
	

	reg PE_add, send_req, send_data_valid;
	reg [7:0] n_ID, src_node, dest_node;

	// unused
	wire unused1;
	wire [63:0] unused2;
	reg [5:0] unused4;
	reg unused5;


	reg [3:0] Node_state;
	localparam START = 4'd0;
	localparam BROADCAST_A = 4'd1;
	localparam DONE = 4'd2;

	//This selects between the add or multiplication PE result for the PE to IF data 
	//wire: 1 sends the add result and 0 sends the mult result
	//assign send_data = PE_add ? PE_add_result : PE_mult_result; 
	//assign send_data = PE_add ? 32'b11111111111111111111111111111111 : 32'b10000000000000000000000000000001; 

	always @ (posedge N_clk) begin
		if(N_rst == 0)
			begin
				Node_state <= START;
				n_ID <= Node_id;
				flit_count <= 4'b0;
		    	src_node <= 8'd7;
				dest_node <= 8'd4;
				send_data_valid <= 1'b0;
				a <= a_in;
				
				
		end

		else 
		  begin
		   //$display("Node%d: a=%b", n_ID, a);
			//$display("The outgoing flit is: %x", if_o_data);
			// send a 2-flit packet from send port 0 to receive port 1
		    
		    vc = 0;
		    PE_add <= 1;
		    //data = 'ha;
		    //if_o_data <= {1'b1 /*valid*/, 1'b1 /*tail*/, dest_node, vc, send_data};
		    if(n_ID == 8'd7)
		      begin
		        case(Node_state)
		          START:
		          begin
		            send_req <= 1'b1;
		            if(req_ack == 1'b1)
		            	begin
		            		Node_state <= BROADCAST_A;
		            		send_req <= 1'b0;
		            	end
		          end
		            
		          BROADCAST_A:
		          begin
		            send_data_valid<=1'b1;
		            if(flit_count == 4'b0)
		            	begin
		            		send_data<=32'b11111111111111111111111111111111;
		            	end
		            else if(flit_count == 4'd1) 
		            	begin
		            		send_data<=32'b10000000000000010000000000000001;
		            	end
		            else 
		            	begin
		            		send_data_valid <= 1'b0;
		            	end

		            
		            
		            flit_count <= flit_count + 1;
		          end
		          
		          DONE:
		          begin
		            
		          end
		          
		        endcase
		      end // end if
		  end // end else
    
		  if((n_ID == 8'd4) && (if_i_flit[72] == 1))
		    begin
		    		$display("Node%d received data is: %b", n_ID, if_i_flit[31:0]);
   		  		 //$display("@%3d: Ejecting flit %x at receive port %0d", cycle, flit_out_wire[i], i);//, nodes[i]);
	      end
		end

	 m_if_2_router_v3 IF_Router(
		.clk(N_clk), .rst_n(N_rst),
		//general sending interface for master pe and mig_office
		//signals between PE and IF
		.i_comm_send_req(send_req),
		.o_comm_send_ack(req_ack),
		.i_data_valid(send_data_valid),
		.i_data(send_data),
		.i_src(src_node),
		.i_dst(dest_node),
		.local_id(n_ID),
		
		
		//signals Between IF and ROUTER
		.i_credit(if_i_credit),
		.o_credit_valid(if_o_credit_valid),
		.o_credit(if_o_credit),
		.o_data(if_o_data),
		.o_data_valid(if_o_data_valid),
		.i_flit(if_i_flit),


		//Unused
		
		.i_id(unused4),
		.i_ack_rx(unused5),
		.o_req_rx(unused1),
		.o_data_input(unused2),
		.o_data_input_valid(unused1),
		.i_seq_len(unused4)
		);


	PE processor_element(.clk(N_clk), .A(test_value_A), .B(test_value_B), 
						.C(test_value_C), .mult_result(PE_mult_result),
						.add_result(PE_add_result));



endmodule



